module hello;

    initial begin
        $display("System Verilog is running");
        $finish;
    end

endmodule